library verilog;
use verilog.vl_types.all;
entity memorysystem is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        nWAIT           : out    vl_logic;
        BIGEND          : out    vl_logic;
        HIVECS          : out    vl_logic;
        ID              : out    vl_logic_vector(31 downto 0);
        IABORT          : out    vl_logic;
        InMREQ          : in     vl_logic;
        InTRANS         : in     vl_logic;
        ISEQ            : in     vl_logic;
        ITBIT           : in     vl_logic;
        IA              : in     vl_logic_vector(31 downto 0);
        InM             : in     vl_logic_vector(4 downto 0);
        DDIN            : out    vl_logic_vector(31 downto 0);
        DABORT          : out    vl_logic;
        DA              : in     vl_logic_vector(31 downto 0);
        DD              : in     vl_logic_vector(31 downto 0);
        DnRW            : in     vl_logic;
        DnMREQ          : in     vl_logic;
        DMAS            : in     vl_logic_vector(1 downto 0);
        DMORE           : in     vl_logic;
        DLOCK           : in     vl_logic;
        DDEN            : in     vl_logic;
        DnTRANS         : in     vl_logic;
        DSEQ            : in     vl_logic;
        DnM             : in     vl_logic_vector(4 downto 0);
        HCLK            : in     vl_logic;
        HRDATAM         : in     vl_logic_vector(31 downto 0);
        HREADYM         : in     vl_logic;
        HRESPM          : in     vl_logic_vector(1 downto 0);
        HGRANTM         : in     vl_logic;
        HADDRM          : out    vl_logic_vector(31 downto 0);
        HTRANSM         : out    vl_logic_vector(1 downto 0);
        HWRITEM         : out    vl_logic;
        HSIZEM          : out    vl_logic_vector(2 downto 0);
        HBURSTM         : out    vl_logic_vector(2 downto 0);
        HPROTM          : out    vl_logic_vector(3 downto 0);
        HWDATAM         : out    vl_logic_vector(31 downto 0);
        HBUSREQM        : out    vl_logic;
        HLOCKM          : out    vl_logic;
        CPID            : in     vl_logic_vector(31 downto 0);
        CPLATECANCEL    : in     vl_logic;
        nCPMREQ         : in     vl_logic;
        CPPASS          : in     vl_logic;
        CPTBIT          : in     vl_logic;
        nCPTRANS        : in     vl_logic;
        CPDOUT          : in     vl_logic_vector(31 downto 0);
        CHSDE           : out    vl_logic_vector(1 downto 0);
        CHSEX           : out    vl_logic_vector(1 downto 0);
        CPEN            : out    vl_logic;
        CPDIN           : out    vl_logic_vector(31 downto 0);
        nfiq            : in     vl_logic;
        nirq            : in     vl_logic;
        CP15protect     : in     vl_logic
    );
end memorysystem;
