library verilog;
use verilog.vl_types.all;
entity Wraper is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        IMMU_HRDATAM    : out    vl_logic_vector(31 downto 0);
        IMMU_HREADYM    : out    vl_logic;
        IMMU_HADDRM     : in     vl_logic_vector(31 downto 0);
        IMMU_HTRANSM    : in     vl_logic_vector(1 downto 0);
        IMMU_HWRITEM    : in     vl_logic;
        IMMU_HSIZEM     : in     vl_logic_vector(2 downto 0);
        IMMU_HBURSTM    : in     vl_logic_vector(2 downto 0);
        IMMU_HPROTM     : in     vl_logic_vector(3 downto 0);
        IMMU_HWDATAM    : in     vl_logic_vector(31 downto 0);
        IMMU_HBUSREQM   : in     vl_logic;
        IMMU_HLOCKM     : in     vl_logic;
        DMMU_HRDATAM    : out    vl_logic_vector(31 downto 0);
        DMMU_HREADYM    : out    vl_logic;
        DMMU_HADDRM     : in     vl_logic_vector(31 downto 0);
        DMMU_HTRANSM    : in     vl_logic_vector(1 downto 0);
        DMMU_HWRITEM    : in     vl_logic;
        DMMU_HSIZEM     : in     vl_logic_vector(2 downto 0);
        DMMU_HBURSTM    : in     vl_logic_vector(2 downto 0);
        DMMU_HPROTM     : in     vl_logic_vector(3 downto 0);
        DMMU_HWDATAM    : in     vl_logic_vector(31 downto 0);
        DMMU_HBUSREQM   : in     vl_logic;
        DMMU_HLOCKM     : in     vl_logic;
        IEXT_HRDATAM    : out    vl_logic_vector(31 downto 0);
        IEXT_HREADYM    : out    vl_logic;
        IEXT_HRESPM     : out    vl_logic_vector(1 downto 0);
        IEXT_HADDRM     : in     vl_logic_vector(31 downto 0);
        IEXT_HTRANSM    : in     vl_logic_vector(1 downto 0);
        IEXT_HWRITEM    : in     vl_logic;
        IEXT_HSIZEM     : in     vl_logic_vector(2 downto 0);
        IEXT_HBURSTM    : in     vl_logic_vector(2 downto 0);
        IEXT_HPROTM     : in     vl_logic_vector(3 downto 0);
        IEXT_HWDATAM    : in     vl_logic_vector(31 downto 0);
        IEXT_HBUSREQM   : in     vl_logic;
        IEXT_HLOCKM     : in     vl_logic;
        DEXT_HRDATAM    : out    vl_logic_vector(31 downto 0);
        DEXT_HREADYM    : out    vl_logic;
        DEXT_HRESPM     : out    vl_logic_vector(1 downto 0);
        DEXT_HADDRM     : in     vl_logic_vector(31 downto 0);
        DEXT_HTRANSM    : in     vl_logic_vector(1 downto 0);
        DEXT_HWRITEM    : in     vl_logic;
        DEXT_HSIZEM     : in     vl_logic_vector(2 downto 0);
        DEXT_HBURSTM    : in     vl_logic_vector(2 downto 0);
        DEXT_HPROTM     : in     vl_logic_vector(3 downto 0);
        DEXT_HWDATAM    : in     vl_logic_vector(31 downto 0);
        DEXT_HBUSREQM   : in     vl_logic;
        DEXT_HLOCKM     : in     vl_logic;
        ICache_HRDATAM  : out    vl_logic_vector(31 downto 0);
        ICache_HREADYM  : out    vl_logic;
        ICache_HADDRM   : in     vl_logic_vector(31 downto 0);
        ICache_HTRANSM  : in     vl_logic_vector(1 downto 0);
        ICache_HWRITEM  : in     vl_logic;
        ICache_HSIZEM   : in     vl_logic_vector(2 downto 0);
        ICache_HBURSTM  : in     vl_logic_vector(2 downto 0);
        ICache_HPROTM   : in     vl_logic_vector(3 downto 0);
        ICache_HWDATAM  : in     vl_logic_vector(31 downto 0);
        ICache_HBUSREQM : in     vl_logic;
        ICache_HLOCKM   : in     vl_logic;
        DCache_HRDATAM  : out    vl_logic_vector(31 downto 0);
        DCache_HREADYM  : out    vl_logic;
        DCache_HADDRM   : in     vl_logic_vector(31 downto 0);
        DCache_HTRANSM  : in     vl_logic_vector(1 downto 0);
        DCache_HWRITEM  : in     vl_logic;
        DCache_HSIZEM   : in     vl_logic_vector(2 downto 0);
        DCache_HBURSTM  : in     vl_logic_vector(2 downto 0);
        DCache_HPROTM   : in     vl_logic_vector(3 downto 0);
        DCache_HWDATAM  : in     vl_logic_vector(31 downto 0);
        DCache_HBUSREQM : in     vl_logic;
        DCache_HLOCKM   : in     vl_logic;
        WB_HRDATAM      : out    vl_logic_vector(31 downto 0);
        WB_HREADYM      : out    vl_logic;
        WB_HADDRM       : in     vl_logic_vector(31 downto 0);
        WB_HTRANSM      : in     vl_logic_vector(1 downto 0);
        WB_HWRITEM      : in     vl_logic;
        WB_HSIZEM       : in     vl_logic_vector(2 downto 0);
        WB_HBURSTM      : in     vl_logic_vector(2 downto 0);
        WB_HPROTM       : in     vl_logic_vector(3 downto 0);
        WB_HWDATAM      : in     vl_logic_vector(31 downto 0);
        WB_HBUSREQM     : in     vl_logic;
        WB_HLOCKM       : in     vl_logic;
        HRDATAM         : in     vl_logic_vector(31 downto 0);
        HREADYM         : in     vl_logic;
        HRESPM          : in     vl_logic_vector(1 downto 0);
        HGRANTM         : in     vl_logic;
        HADDRM          : out    vl_logic_vector(31 downto 0);
        HTRANSM         : out    vl_logic_vector(1 downto 0);
        HWRITEM         : out    vl_logic;
        HSIZEM          : out    vl_logic_vector(2 downto 0);
        HBURSTM         : out    vl_logic_vector(2 downto 0);
        HPROTM          : out    vl_logic_vector(3 downto 0);
        HWDATAM         : out    vl_logic_vector(31 downto 0);
        HBUSREQM        : out    vl_logic;
        HLOCKM          : out    vl_logic
    );
end Wraper;
