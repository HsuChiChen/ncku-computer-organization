library verilog;
use verilog.vl_types.all;
entity Direct_Map_D_Cache is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        nWAIT           : in     vl_logic;
        BIGEND          : in     vl_logic;
        Invalid_DCache  : in     vl_logic;
        Invalid_DCache_MVA: in     vl_logic;
        Clean_DCache_MVA: in     vl_logic;
        Clean_Invalid_DCache_MVA: in     vl_logic;
        Clean_DCache_Index: in     vl_logic;
        Clean_Invalid_DCache_Index: in     vl_logic;
        Entry_MVA_Index : in     vl_logic_vector(26 downto 0);
        Data_phase_Cacheable: in     vl_logic;
        Data_phase_Bufferable: in     vl_logic;
        nMREQ           : in     vl_logic;
        MVA             : in     vl_logic_vector(31 downto 0);
        Data_phase_MAS  : in     vl_logic_vector(1 downto 0);
        Data_phase_nRW  : in     vl_logic;
        DO              : in     vl_logic_vector(31 downto 0);
        DI              : out    vl_logic_vector(31 downto 0);
        Cache_nWAIT     : out    vl_logic;
        fill            : out    vl_logic;
        Data_phase_MVA  : in     vl_logic_vector(31 downto 0);
        fill_finish     : in     vl_logic;
        TAG_WAddr       : in     vl_logic_vector(26 downto 0);
        TAG_WE          : in     vl_logic;
        Valid_WAddr     : in     vl_logic_vector(1 downto 0);
        Valid_WE        : in     vl_logic;
        Valid_WData     : in     vl_logic;
        Value_WAddr     : in     vl_logic_vector(4 downto 0);
        Value_WE        : in     vl_logic_vector(3 downto 0);
        Value_WData     : in     vl_logic_vector(31 downto 0);
        PA_TAG_WAddr    : in     vl_logic_vector(1 downto 0);
        PA_TAG_WE       : in     vl_logic;
        PA_TAG_WData    : in     vl_logic_vector(25 downto 0);
        Dirty_WAddr     : in     vl_logic_vector(1 downto 0);
        Dirty_WE        : in     vl_logic_vector(1 downto 0);
        Dirty_WData     : in     vl_logic_vector(1 downto 0);
        Retry           : out    vl_logic;
        Data_phase_Cache_Hit: out    vl_logic;
        Cache_operation_EN: out    vl_logic;
        Write_Back      : out    vl_logic;
        Write_Back_Addr : out    vl_logic_vector(27 downto 0);
        Write_Back_Data : out    vl_logic_vector(127 downto 0);
        Write_Back_nWAIT: in     vl_logic
    );
end Direct_Map_D_Cache;
