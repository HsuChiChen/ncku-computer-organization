`timescale 10ns / 1ps

module testbench;

	reg		[31:0]	ins;
	
	wire	[31:0]	op1, op2;
	wire	[3:0]	aluop;
	
	DECODE decode (op1, op2, aluop, ins);
	
	initial
	begin
		// zero
		ins = 32'b00000000000000000000000000000000;
		#100;
		// ADD	a5,a2,a3  aluop=0000  op1=24  op2=26
		ins = 32'b00000000110101100000011110110011;
		#100;
		// ADDI	a5,a2,15  aluop=0000  op1=24  op2=15
		ins = 32'b00000000111101100000011110010011;
		#100;
		// SUB	a5,a2,a3  aluop=1000  op1=24  op2=26
		ins = 32'b01000000110101100000011110110011;
		#100;
		// AND	a5,a2,a3  aluop=0111  op1=24  op2=26
		ins = 32'b00000000110101100111011110110011;
		#100;
		// ANDI	a5,a2,4   aluop=0111  op1=24  op2=4
		ins = 32'b00000000010001100111011110010011;
		#100;
		// OR	a5,a2,a3  aluop=0110  op1=24  op2=26
		ins = 32'b00000000110101100110011110110011;
		#100;
		// ORI	a5,a2,2   aluop=0110  op1=24  op2=2
		ins = 32'b00000000001001100110011110010011;
		#100;
		// XOR	a5,a2,a3  aluop=0100  op1=24  op2=26
		ins = 32'b00000000110101100100011110110011;
		#100;
		// XORI	a5,a2,1   aluop=0100  op1=24  op2=1
		ins = 32'b00000000000101100100011110010011;
		#100;
		// SLT	a5,a3,a2  aluop=0010  op1=26  op2=24
		ins = 32'b00000000110001101010011110110011;
		#100;
		// SLTI	a5,a3,4   aluop=0010  op1=26  op2=4
		ins = 32'b00000000010001101010011110010011;
		#100;
		// SLTU	a5,a4,a2  aluop=0011  op1=28  op2=24
		ins = 32'b00000000110001110011011110110011;
		#100;
		// SLTIU a5,a3,8  aluop=0011  op1=26  op2=8
		ins = 32'b00000000100001101011011110010011;
		#100;
		// SLL	a5,a3,a2  aluop=0001  op1=26  op2=24
		ins = 32'b00000000110001101001011110110011;
		#100;
		// SRL	a5,a3,a2  aluop=0101  op1=26  op2=24
		ins = 32'b00000000110001101101011110110011;
		#100;
		// SRA	a5,a4,a2  aluop=1101  op1=28  op2=24
		ins = 32'b01000000110001110101011110110011;
		#200 $stop;
	end
endmodule
		