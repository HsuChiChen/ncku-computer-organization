library verilog;
use verilog.vl_types.all;
entity exe_bypassing is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        nWAIT           : in     vl_logic;
        load_pc_flush   : in     vl_logic;
        cause_exception : in     vl_logic;
        updated_cpsr    : in     vl_logic_vector(31 downto 0);
        id_exe_write_addr: in     vl_logic_vector(3 downto 0);
        id_mem_write_addr: in     vl_logic_vector(3 downto 0);
        ctl_load_data_width: in     vl_logic_vector(1 downto 0);
        ctl_load_data_sign: in     vl_logic;
        swap_enable     : in     vl_logic;
        chk_branch      : in     vl_logic;
        chk_exe_write_enable: in     vl_logic;
        chk_mem_write_enable: in     vl_logic;
        chk_branch_link : in     vl_logic;
        ctl_multiply_type: in     vl_logic_vector(2 downto 0);
        ctl_psr_write_mask: in     vl_logic_vector(3 downto 0);
        chk_psr_write_enable: in     vl_logic;
        ctl_psr_sel     : in     vl_logic;
        ctl_data_from_mem: in     vl_logic;
        back_from_exception: in     vl_logic;
        ctl_lw_str_instruction: in     vl_logic;
        exe_swap_enable : out    vl_logic;
        exe_write_addr  : out    vl_logic_vector(3 downto 0);
        exe_bypass_write_enable: out    vl_logic;
        exe_mem_write_addr: out    vl_logic_vector(3 downto 0);
        exe_mem_write_enable: out    vl_logic;
        exe_load_data_width: out    vl_logic_vector(1 downto 0);
        exe_load_data_sign: out    vl_logic;
        exe_multiply_type: out    vl_logic_vector(2 downto 0);
        exe_data_from_mem: out    vl_logic;
        exe_psr_write_mask: out    vl_logic_vector(3 downto 0);
        exe_psr_write_enable: out    vl_logic;
        exe_psr_write_data: out    vl_logic_vector(31 downto 0);
        exe_psr_sel     : out    vl_logic;
        back_to_usr_mode: out    vl_logic;
        exe_branch_link : out    vl_logic;
        exe_branch      : out    vl_logic;
        exe_lw_str_instruction: out    vl_logic;
        ctl_mrs_instruction: in     vl_logic;
        exe_mrs_instruction: out    vl_logic;
        ldm2            : in     vl_logic;
        exe_ldm2        : out    vl_logic
    );
end exe_bypassing;
