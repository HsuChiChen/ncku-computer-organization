library verilog;
use verilog.vl_types.all;
entity TBTic is
    generic(
        PERIOD          : integer := 10
    );
end TBTic;
