library verilog;
use verilog.vl_types.all;
entity EASY is
    port(
        HCLK            : in     vl_logic;
        HRESETn         : in     vl_logic
    );
end EASY;
