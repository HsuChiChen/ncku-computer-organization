
module DECODE (op1, op2, aluop, ins);

	input 	[31:0]	ins;

    output  [31:0]  op1;
    output  [31:0]  op2;
    output  [3:0]   aluop;

	wire	[6:0]	opcode, funct7;
	wire	[4:0]	rs1, rs2, rd;
	wire    [2:0]   funct3;
    reg     [31:0]  REG [0:32];
    integer i;
    
    // initial REG data  
    initial begin
        for(i = 0; i < 32; i = i + 1) begin
            REG[i] = i*2;
        end
    end

    //=======================================================================
    // R-type
    // | 31      25 | 24   20 | 19   15 | 14      12 | 11  07 | 06      00 |
    // +------------+---------+---------+------------+--------+------------+
    // |   funct7   |   rs2   |   rs1   |   funct3   |   rd   |   opcode   |
    // +------------+---------+---------+------------+--------+------------+
    //     0000000       add                000                   0110011
    //     0100000       sub                000                   0110011
    //     0000000       shl                001                   0110011
    //     0000000       slt                010                   0110011
    //     0000000       sltu               011                   0110011 
    //     0000000       xor                100                   0110011 
    //     0000000       shr                101                   0110011
    //     0100000       shra               101                   0110011
    //     0000000       or                 110                   0110011 
    //     0000000       and                111                   0110011 
    //
    // ---------------------------------------------------------------------
    // I-type
    // | 31                20 | 19   15 | 14      12 | 11  07 | 06      00 |
    // +----------------------+---------+------------+--------+------------+
    // |   immediate[11:0]    |   rs1   |   funct3   |   rd   |   opcode   |
    // +----------------------+---------+------------+--------+------------+
    //            addi                       000                  0010011
    //            slti                       010                  0010011
    //            sltiu                      011                  0010011
    //            xori                       100                  0010011
    //            ori                        110                  0010011
    //            andi                       111                  0010011
    //
    //=======================================================================

    assign opcode = ins[6:0];
    assign rs1 = ins[19:15];
    assign rs2 = (opcode[6:0] == 7'b0110011)?ins[24:20]:5'd0;
    assign rd  = ins[11:7];
    assign funct3 = ins[14:12];
    assign funct7 = (opcode[6:0] == 7'b0110011)?ins[31:25]:7'd0;

    assign op1 = REG[rs1];
    assign op2 = (opcode[6:0] == 7'b0110011)?REG[rs2]:ins[31:20];

    //=============================================
    // Ins   		funct7      funct3     ALUOP	
    // +-----------+----------+----------+--------+
    // ADD	        0000000     000        0000	
    // ADDI         -           000        0000
    // SUB		    0100000     000        1000	
    // SLT		    0000000     010        0010	
    // SLTI         -           010        0010
    // SLTU	        0000000     011        0011
    // SLTIU        -           011        0011
    // XOR		    0000000     100        0100	
    // XORI         -           100        0100
    // OR		    0000000     110        0110	
    // ORI          -           110        0110
    // AND          0000000     111        0111
    // ANDI         -           111        0111
    // SLL		    0000000     001        0001	
    // SRL		    0000000     101        0101	
    // SRA	        0100000     101        1101	
    //=============================================

    assign aluop = (opcode[6:0] == 7'b0110011)?{funct7[5], funct3}:{1'b0, funct3};

endmodule