module reg00
(
    input  logic [31:0] x0,
    input  logic [31:0] x1,
    input  logic [31:0] x2,
    input  logic [31:0] x3,
    input  logic [31:0] x4,
    input  logic [31:0] x5,
    input  logic [31:0] x6,
    input  logic [31:0] x7,
    input  logic [31:0] x8,
    input  logic [31:0] x9,
    input  logic [31:0] x10,
    input  logic [31:0] x11,
    input  logic [31:0] x12,
    input  logic [31:0] x13,
    input  logic [31:0] x14,
    input  logic [31:0] x15,
    input  logic [31:0] x16,
    input  logic [31:0] x17,
    input  logic [31:0] x18,
    input  logic [31:0] x19,
    input  logic [31:0] x20,
    input  logic [31:0] x21,
    input  logic [31:0] x22,
    input  logic [31:0] x23,
    input  logic [31:0] x24,
    input  logic [31:0] x25,
    input  logic [31:0] x26,
    input  logic [31:0] x27,
    input  logic [31:0] x28,
    input  logic [31:0] x29,
    input  logic [31:0] x30,
    input  logic [31:0] x31

);

endmodule
