library verilog;
use verilog.vl_types.all;
entity WFI is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        nWAIT           : in     vl_logic;
        Wait_for_interrupt: in     vl_logic;
        nfiq            : in     vl_logic;
        nirq            : in     vl_logic;
        WFI_nWAIT       : out    vl_logic
    );
end WFI;
