library verilog;
use verilog.vl_types.all;
entity general_regs is
    port(
        clk             : in     vl_logic;
        rst_n           : in     vl_logic;
        nWAIT           : in     vl_logic;
        HIVECS          : in     vl_logic;
        load_pc_flush   : in     vl_logic;
        stall_instruction_fetch: in     vl_logic;
        immed_value_sel : in     vl_logic_vector(2 downto 0);
        fourth_addr_sel : in     vl_logic_vector(1 downto 0);
        multiple_store  : in     vl_logic;
        str_instruction : in     vl_logic;
        multiply_mula   : in     vl_logic;
        swap_enable     : in     vl_logic;
        chk_branch      : in     vl_logic;
        ctl_branch_link : in     vl_logic;
        exe_branch_link : in     vl_logic;
        mem_write_enable: in     vl_logic;
        mem_write_addr  : in     vl_logic_vector(3 downto 0);
        mem_write_data  : in     vl_logic_vector(31 downto 0);
        exe_write_enable: in     vl_logic;
        exe_write_addr  : in     vl_logic_vector(3 downto 0);
        exe_write_data  : in     vl_logic_vector(31 downto 0);
        ctl_lw_str_instruction: in     vl_logic;
        multiple_finished: in     vl_logic;
        multiple_last   : in     vl_logic;
        data_abort      : in     vl_logic;
        cause_exception : in     vl_logic;
        what_exception  : in     vl_logic_vector(2 downto 0);
        back_to_usr_mode: in     vl_logic;
        write_to_regpc  : in     vl_logic_vector(31 downto 0);
        return_addr     : in     vl_logic_vector(31 downto 0);
        fet_condition_code: in     vl_logic_vector(3 downto 0);
        psr_mode        : in     vl_logic_vector(4 downto 0);
        id_first_opern  : out    vl_logic_vector(31 downto 0);
        id_second_opern : out    vl_logic_vector(31 downto 0);
        id_third_opern  : out    vl_logic_vector(31 downto 0);
        id_fourth_opern : out    vl_logic_vector(31 downto 0);
        id_regpc        : out    vl_logic_vector(31 downto 0);
        id_first_addr   : out    vl_logic_vector(3 downto 0);
        id_second_addr  : out    vl_logic_vector(3 downto 0);
        id_third_addr   : out    vl_logic_vector(3 downto 0);
        id_fourth_addr  : out    vl_logic_vector(3 downto 0);
        id_condition_code: out    vl_logic_vector(3 downto 0);
        id_exe_write_addr: out    vl_logic_vector(3 downto 0);
        id_mem_write_addr: out    vl_logic_vector(3 downto 0);
        immed_value     : out    vl_logic_vector(31 downto 0);
        instruction     : in     vl_logic_vector(31 downto 0);
        mem_lw_str_instruction: in     vl_logic;
        multiple_end    : in     vl_logic;
        Fourth_ADDR     : out    vl_logic_vector(3 downto 0);
        stm2            : in     vl_logic;
        mem_ldm2        : in     vl_logic;
        stall_delay     : in     vl_logic
    );
end general_regs;
